entity mux is
    port (
        clk: in std_logic
    );
end entity mux;