entity ctrl_unit is
    port (
        clk: in std_logic;
    );
end entity ctrl_unit;