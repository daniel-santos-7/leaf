package body core_pkg is
    
    constant word_size: natural := 32;

    constant instruction_size: natural := 32;
    
end package body core_pkg;