entity branch_predictor is
    port (
        clk: in std_logic
    );
end entity branch_predictor;