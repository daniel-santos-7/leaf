entity demux is
    port (
        clk: in std_logic;
    );
end entity demux;